module tlk2711_tb();


endmodule