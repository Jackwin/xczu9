module top (

input       sys_clk_50,
input       sys_rstn

);

endmodule