
///////////////////////////////////////////////////////////////////////////////
//  
//    Version: 1.0
//    Filename:  tlk2711_top.v
//    Date Created: 2021-06-27
// 
//   
// Project: TLK2711
// Device: zu9eg
// Purpose: top file
// Author: Zhu Lin
// Reference:  
// Revision History:
//   Rev 1.0 - First created, zhulin, 2021-07-03
//   
// Email: 
////////////////////////////////////////////////////////////////////////////////

module tlk2711_top 
#(       
    parameter DEBUG_ENA = "TRUE",
    parameter ADDR_WIDTH = 48,
    parameter AXI_RDATA_WIDTH = 64,
    parameter AXI_WDATA_WIDTH = 64,
    parameter AXI_WBYTE_WIDTH = 8,
    parameter STREAM_RDATA_WIDTH = 64,
    parameter STREAM_WDATA_WIDTH = 64,
    parameter STREAM_WBYTE_WIDTH = 8,
    parameter DLEN_WIDTH = 16,

    parameter ADDR_MASK = 16'h00ff,
    parameter ADDR_BASE = 16'h0000
)
(  
    input               ps_clk,
    input               ps_rst,
    
    //register config
    input               i_reg_wen,
    input  [15:0]       i_reg_waddr,
    input  [63:0]       i_reg_wdata,
    
    //register status 
    input               i_reg_ren,
    input  [15:0]       i_reg_raddr,
    output [63:0]       o_reg_rdata,
    
    //interrupt
    output              o_tx_irq,
    output              o_rx_irq,
    output              o_loss_irq,

    //tlk2711 interface
    input               clk,
    input               rst,

    input               i_2711_rkmsb,
    input               i_2711_rklsb,
    input   [15:0]      i_2711_rxd,
    output              o_2711_tkmsb,
    output              o_2711_tklsb,
    output              o_2711_enable,
    output              o_2711_loopen,
    output              o_2711_lckrefn,
    output              o_2711_testen,
    output              o_2711_prbsen,
    output              o_2711_pre,
    output  [15:0]      o_2711_txd,

    //PS interface  
    //AXI4 Memory Mapped Read Address Interface Signals
    input           m_axi_arready,
    output          m_axi_arvalid,
    output [3:0]    m_axi_arid,
    output [ADDR_WIDTH-1:0] m_axi_araddr,
    output [7:0]    m_axi_arlen,
    output [2:0]    m_axi_arsize,
    output [1:0]    m_axi_arburst,
    output [2:0]    m_axi_arprot,
    output [3:0]    m_axi_arcache,
    output          m_axi_aruser,
   
    //AXI4 Memory Mapped Read Data Interface Signals
    input [AXI_RDATA_WIDTH-1:0]   m_axi_rdata,
    input [1:0]     m_axi_rresp,
    input           m_axi_rlast,
    input           m_axi_rvalid,
    output          m_axi_rready,

    //AXI4 Memory Mapped Write Address Interface Signals
    input           m_axi_awready,
    output          m_axi_awvalid,
    output [3:0]    m_axi_awid,
    output [ADDR_WIDTH-1:0]   m_axi_awaddr,
    output [7:0]    m_axi_awlen,
    output [2:0]    m_axi_awsize,
    output [1:0]    m_axi_awburst,
    output [2:0]    m_axi_awprot,
    output [3:0]    m_axi_awcache,
    output [3:0]    m_axi_awuser,   

    //AXI4 Memory Mapped Write Data Interface Signals
    output [AXI_WDATA_WIDTH-1:0]  m_axi_wdata,
    output [AXI_WBYTE_WIDTH-1:0]  m_axi_wstrb,
    output          m_axi_wlast,
    output          m_axi_wvalid,
    input           m_axi_wready,

    input [1:0]     m_axi_bresp,
    input           m_axi_bvalid,
    output          m_axi_bready
   
);

    wire [ADDR_WIDTH-1:0]   tx_base_addr;
    wire [31:0]             tx_total_length;
    wire [15:0]             tx_packet_body;
    wire [15:0]             tx_packet_tail;
    wire [23:0]             tx_body_num;
    wire [2:0]              tx_mode;
    wire                    loopback_ena;
    wire                    tx_config_done; 
    wire                    tx_interrupt;
    wire                    tx_pre;

    wire [ADDR_WIDTH-1:0]   rx_base_addr;
    wire                    rx_config_done;
    wire                    rx_interrupt;
    wire [15:0]             rx_frame_length;
    wire [15:0]             rx_packet_body; 
    wire [15:0]             rx_packet_tail;
    wire [23:0]             rx_frame_num;
    wire [23:0]             line_num_per_intr;
    wire [19:0]             backward_cycle_num;

    wire [15:0]             tx_intr_width;
    wire [15:0]             rx_intr_width;
    wire [15:0]             link_intr_width;

    wire                    loss_interrupt;
    wire                    sync_loss;
    wire                    link_loss;
    wire                    soft_rst;
    wire [3:0]              rx_data_type;
    wire                    rx_file_end_flag;
    wire                    rx_checksum_flag;
    wire [1:0]              rx_channel_id;

    wire [DLEN_WIDTH+ADDR_WIDTH-1:0]    rd_cmd_data;
    wire                                rd_cmd_req;
    wire                                rd_cmd_ack;
    wire [DLEN_WIDTH+ADDR_WIDTH-1:0]    wr_cmd_data;
    wire                                wr_cmd_req;
    wire                                wr_cmd_ack;

    wire                                dma_rd_ready;
    wire                                dma_rd_valid;
    wire                                dma_rd_last;
    wire [STREAM_RDATA_WIDTH-1:0]       dma_rd_data;

    wire                                dma_wr_valid;
    wire [STREAM_WBYTE_WIDTH-1:0]       dma_wr_keep;
    wire [STREAM_WDATA_WIDTH-1:0]       dma_wr_data;
    wire                                dma_wr_ready;
    wire                                wr_finish;
            
    wire [10:0]                         rx_status;
    wire [9:0]                          tx_status;
    wire                                rx_fifo_rd;
    wire                                link_loss_detect_ena;
    wire                                sync_loss_detect_ena;
    wire                                check_ena;
    wire                                rx_length_unit;
    wire                                tx_stop_test;
    //wire                                rx_start_test;
    wire [3:0]                          rx_test_error;

   reg_mgt #(
       .DEBUG_ENA(DEBUG_ENA),
       .ADDR_WIDTH(ADDR_WIDTH),
       .ADDR_MASK(ADDR_MASK),
       .ADDR_BASE(ADDR_BASE)
   ) reg_mgt (  
       .ps_clk(ps_clk),
       .ps_rst(ps_rst),
       .i_reg_wen(i_reg_wen),
       .i_reg_waddr(i_reg_waddr),
       .i_reg_wdata(i_reg_wdata),
       .i_reg_ren(i_reg_ren),
       .i_reg_raddr(i_reg_raddr),
       .o_reg_rdata(o_reg_rdata),
       .o_tx_irq(o_tx_irq),
       .o_rx_irq(o_rx_irq),
       .o_loss_irq(o_loss_irq),
       .o_tx_intr_width(tx_intr_width),
       .o_rx_intr_width(rx_intr_width),
       .o_link_intr_width(link_intr_width),

       .clk(clk),
       .rst(rst),
       .o_tx_base_addr(tx_base_addr), 
       .o_tx_total_length(tx_total_length), 
       .o_tx_packet_body(tx_packet_body), 
       .o_tx_packet_tail(tx_packet_tail), 
       .o_tx_body_num(tx_body_num),  
       .o_tx_mode(tx_mode), 
       .o_loopback_ena(loopback_ena),
       .o_tx_config_done(tx_config_done),
       .o_tx_stop_test(tx_stop_test),
       .i_tx_interrupt(tx_interrupt), 
       .o_tx_pre(tx_pre),
       .o_line_num_per_intr(line_num_per_intr),
       .o_backward_cycle_num(backward_cycle_num),

       .o_rx_base_addr(rx_base_addr), 
       .o_rx_config_done(rx_config_done),
      // .o_rx_start_test(rx_start_test),
       .o_rx_fifo_rd(rx_fifo_rd),
       .o_link_loss_detect_ena(link_loss_detect_ena),
       .o_sync_loss_detect_ena(sync_loss_detect_ena),
       .o_rx_check_ena(check_ena),
       .o_rx_length_unit(rx_length_unit),

       .i_rx_interrupt(rx_interrupt), 
       .i_rx_frame_length(rx_frame_length),
       .i_rx_frame_num(rx_frame_num),
       .i_rx_data_type(rx_data_type),
       .i_rx_file_end_flag(rx_file_end_flag),
       .i_rx_checksum_flag(rx_checksum_flag),
       .i_rx_channel_id(rx_channel_id),
      // .i_rx_test_check_error(rx_test_check_error),
       //.i_rx_test_error_status(rx_test_error_status),
       
       .i_tx_status(tx_status),
       .i_rx_test_error(rx_test_error),
       .i_rx_status(rx_status),
       .i_loss_interrupt(loss_interrupt),
       .i_sync_loss(sync_loss),
       .i_link_loss(link_loss),
       .o_soft_rst(soft_rst) 
    );
 
    tlk2711_dma #(
        .AXI_RDATA_WIDTH(AXI_RDATA_WIDTH),
        .AXI_WDATA_WIDTH(AXI_WDATA_WIDTH), 
        .AXI_WBYTE_WIDTH(AXI_WBYTE_WIDTH), 
        .STREAM_RDATA_WIDTH(STREAM_RDATA_WIDTH),
        .STREAM_WDATA_WIDTH(STREAM_WDATA_WIDTH), 
        .STREAM_WBYTE_WIDTH(STREAM_WBYTE_WIDTH),   
        .ADDR_WIDTH(ADDR_WIDTH),
        .DLEN_WIDTH(DLEN_WIDTH)  
    ) tlk2711_dma (
        .clk(clk),
        .rst(rst),
        .i_rd_cmd_data(rd_cmd_data), 
        .i_rd_cmd_req(rd_cmd_req),
        .o_rd_cmd_ack(rd_cmd_ack),
        .i_wr_cmd_data(wr_cmd_data), 
        .i_wr_cmd_req(wr_cmd_req),
        .o_wr_cmd_ack(wr_cmd_ack),
        .i_dma_rd_ready(dma_rd_ready),
        .o_dma_rd_valid(dma_rd_valid),
        .o_dma_rd_last(dma_rd_last),
        .o_dma_rd_data(dma_rd_data),
        .i_dma_wr_valid(dma_wr_valid),
        .i_dma_wr_keep(dma_wr_keep),
        .i_dma_wr_data(dma_wr_data),
        .o_dma_wr_ready(dma_wr_ready),
        .o_wr_finish(wr_finish),
        .m_axi_arready(m_axi_arready),
        .m_axi_arvalid(m_axi_arvalid),
        .m_axi_arid(m_axi_arid),
        .m_axi_araddr(m_axi_araddr),
        .m_axi_arlen(m_axi_arlen),
        .m_axi_arsize(m_axi_arsize),
        .m_axi_arburst(m_axi_arburst),
        .m_axi_arprot(m_axi_arprot),
        .m_axi_arcache(m_axi_arcache),
        .m_axi_aruser(m_axi_aruser),
        .m_axi_rdata(m_axi_rdata),
        .m_axi_rresp(m_axi_rresp),
        .m_axi_rlast(m_axi_rlast),
        .m_axi_rvalid(m_axi_rvalid),
        .m_axi_rready(m_axi_rready),
        .m_axi_awready(m_axi_awready),
        .m_axi_awvalid(m_axi_awvalid),
        .m_axi_awid(m_axi_awid),
        .m_axi_awaddr(m_axi_awaddr),
        .m_axi_awlen(m_axi_awlen),
        .m_axi_awsize(m_axi_awsize),
        .m_axi_awburst(m_axi_awburst),
        .m_axi_awprot(m_axi_awprot),
        .m_axi_awcache(m_axi_awcache),
        .m_axi_awuser(m_axi_awuser),   
        .m_axi_wdata(m_axi_wdata),
        .m_axi_wstrb(m_axi_wstrb),
        .m_axi_wlast(m_axi_wlast),
        .m_axi_wvalid(m_axi_wvalid),
        .m_axi_wready(m_axi_wready),
        .m_axi_bresp(m_axi_bresp),
        .m_axi_bvalid(m_axi_bvalid),
        .m_axi_bready(m_axi_bready)
    );

    // reg         tx_start;
    // reg [2:0]   tx_cfg_done;
    // reg [2:0]   rx_cfg_done;
    // reg         rx_start;

    // always @(posedge clk) begin
    //     tx_cfg_done <= {tx_cfg_done[1:0], tx_config_done};
    //     rx_cfg_done <= {rx_cfg_done[1:0], rx_config_done};
    //     tx_start <= ~tx_cfg_done[2] & tx_cfg_done[1];
    //     rx_start <= ~rx_cfg_done[2] & rx_cfg_done[1];
    // end

    tlk2711_tx_cmd #(
        .DEBUG_ENA(DEBUG_ENA),
        .ADDR_WIDTH(ADDR_WIDTH),
        .DLEN_WIDTH(DLEN_WIDTH) 
    ) tlk2711_tx_cmd (
        .clk(clk),
        .rst(rst),
        .i_soft_rst(soft_rst),
        .i_rd_cmd_ack(rd_cmd_ack),
        .o_rd_cmd_req(rd_cmd_req),
        .o_rd_cmd_data(rd_cmd_data), 
        .i_dma_rd_last(dma_rd_last),
        .i_tx_mode(tx_mode), 
        .i_tx_start(tx_config_done),
        .i_tx_base_addr(tx_base_addr),
        .i_tx_packet_body(tx_packet_body), 
        .i_tx_packet_tail(tx_packet_tail), 
        .i_tx_body_num(tx_body_num)
    );

    tlk2711_tx_data #(
        .DEBUG_ENA(DEBUG_ENA),
        .DATA_WIDTH(STREAM_RDATA_WIDTH)
    ) tlk2711_tx_data (
        .clk(clk),
        .rst(rst),
        .i_soft_reset(soft_rst),
        .i_stop_test(tx_stop_test),
        .i_tx_mode(tx_mode),
        .i_loopback_ena(loopback_ena),
        .i_tx_start(tx_config_done),
        .i_tx_packet_body(tx_packet_body), 
        .i_tx_packet_tail(tx_packet_tail),
        .i_tx_body_num(tx_body_num),
        .i_tx_intr_width(tx_intr_width),
        .i_backward_cycle_num(backward_cycle_num),
        .i_tx_pre(tx_pre),
        .i_dma_rd_valid(dma_rd_valid),
        .i_dma_rd_last(dma_rd_last),
        .i_dma_rd_data(dma_rd_data),
        .o_dma_rd_ready(dma_rd_ready),
        .o_tx_interrupt(tx_interrupt),
        .o_tx_status(tx_status),
        .o_2711_tkmsb(o_2711_tkmsb),
        .o_2711_tklsb(o_2711_tklsb),
        .o_2711_enable(o_2711_enable),
        .o_2711_loopen(o_2711_loopen),
        .o_2711_lckrefn(o_2711_lckrefn),
        .o_2711_testen(o_2711_testen),
        .o_2711_prbsen(o_2711_prbsen),
        .o_2711_pre(o_2711_pre),
        .o_2711_txd(o_2711_txd)
    );

    tlk2711_rx_link #(
        .DEBUG_ENA(DEBUG_ENA),
        .ADDR_WIDTH(ADDR_WIDTH),
        .DLEN_WIDTH(DLEN_WIDTH), 
        .DATA_WIDTH(STREAM_RDATA_WIDTH),
        .WBYTE_WIDTH(STREAM_WBYTE_WIDTH)
    ) tlk2711_rx_link (
        .clk(clk),
        .rst(rst),
        .i_soft_rst(soft_rst),
        //.i_rx_start_test(rx_start_test),
        .i_tx_mode(tx_mode), 
        .i_wr_cmd_ack(wr_cmd_ack),
        .o_wr_cmd_req(wr_cmd_req),
        .o_wr_cmd_data(wr_cmd_data), 
        .i_rx_start(rx_config_done),
        .i_rx_base_addr(rx_base_addr),
        .i_rx_line_num_per_intr(line_num_per_intr),
        .i_rx_intr_width(rx_intr_width),
        .i_link_intr_width(link_intr_width),
        .i_link_loss_detect_ena(link_loss_detect_ena),
        .i_sync_loss_detect_ena(sync_loss_detect_ena),
        .i_check_ena(check_ena),
        .i_rx_length_unit(rx_length_unit),
        .i_rx_fifo_rd(rx_fifo_rd),
        .i_dma_wr_ready(dma_wr_ready),
        .i_wr_finish(wr_finish),
        .o_dma_wr_valid(dma_wr_valid),
        .o_dma_wr_keep(dma_wr_keep),
        .o_dma_wr_data(dma_wr_data),
        .o_rx_interrupt(rx_interrupt),
        .o_rx_frame_length(rx_frame_length),
        .o_rx_frame_num(rx_frame_num),
        .o_rx_data_type(rx_data_type),
        .o_rx_file_end_flag(rx_file_end_flag),
        .o_rx_checksum_flag(rx_checksum_flag),
        .o_rx_channel_id(rx_channel_id),
        
        .i_2711_rkmsb(i_2711_rkmsb),
        .i_2711_rklsb(i_2711_rklsb),
        .i_2711_rxd(i_2711_rxd),
        .o_rx_status(rx_status),
        .o_rx_test_error(rx_test_error),
        .o_loss_interrupt(loss_interrupt),
        .o_sync_loss(sync_loss),
        .o_link_loss(link_loss)
    );

    

endmodule

    

    




